always @ (inc,cnt)     //next_cnt 
