`timescale 1ns /1ns

module register16_tb();

